-- part of the solution of exercise 11, chapter 4

package int_package is
    type int_set is array(integer range <>) of integer;
end package int_package;
